* C:\Users\jcasa\Documents\projects\Disruptocooler\pspice\generator.sch

* Schematics Version 9.1 - Web Update 1
* Fri Sep 26 09:25:39 2014



** Analysis setup **
.tran 0ns 5us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "C:\Users\jcasa\Documents\projects\Disruptocooler\pspice\IR2110.sub"
.lib "nom.lib"

.INC "generator.net"
.INC "generator.als"


.probe


.END
